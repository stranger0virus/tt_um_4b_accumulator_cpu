`default_nettype none
`timescale 1ns / 1ps

/* This testbench just instantiates the module and makes some convenient wires
   that can be driven / tested by the cocotb test.py.
*/
module tb ();

  // Dump the signals to a FST file. You can view it with gtkwave or surfer.
  initial begin
    $dumpfile("tb.fst");
    $dumpvars(0, tb);
    #1;
  end

  // Wire up the inputs and outputs:
  reg clk;
  reg rst_n;
  reg ena;
  reg [7:0] ui_in;
  reg [7:0] uio_in;
  wire [7:0] uo_out;
  wire [7:0] uio_out;
  wire [7:0] uio_oe;
`ifdef GL_TEST
  wire VPWR = 1'b1;
  wire VGND = 1'b0;
`endif

  // Replace tt_um_example with your module name:
  tt_um_4b_tiny_cpu user_project (

      // Include power ports for the Gate Level test:
`ifdef GL_TEST
      .VPWR(VPWR),
      .VGND(VGND),
`endif

      .ui_in  (ui_in),    // Dedicated inputs
      .uo_out (uo_out),   // Dedicated outputs
      .uio_in (uio_in),   // IOs: Input path
      .uio_out(uio_out),  // IOs: Output path
      .uio_oe (uio_oe),   // IOs: Enable path (active high: 0=input, 1=output)
      .ena    (ena),      // enable - goes high when design is selected
      .clk    (clk),      // clock
      .rst_n  (rst_n)     // not reset
  );

/*    initial begin

    $monitor("Time=%0t | Input = %b | Sel = %b | Output = %b |  | Imm = %b", $time, ui_in, uio_in, uo_out, uut.imm);
    
	clk   = 0;
    rst_n = 0;
    ui_in = 8'h00;
	uio_in = 8'h00;

    #10 rst_n = 1;
	#5;
	
	ui_in = 8'b00100001;
	uio_in = 8'b00000000;
	#10;

	ui_in = 8'b00110001;
	uio_in = 8'b00000000;
	#10;

    ui_in = 8'b01000010;
    uio_in = 8'b00000000;
    #10;

    ui_in = 8'b01010010;
    uio_in = 8'b00000000;
    #10;

	ui_in = 8'b00100001;
	uio_in = 8'b00000001;
	#300;
        
        $finish;
    end
*/
endmodule
   
